module character_sprites(input [7:0]	addr,
			 output [31:0]	data
			);

	parameter ADDR_WIDTH = 8;
   	parameter DATA_WIDTH =  32;

	// ROM definition
	parameter [0:159][31:0] ROM = {
	
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00011111001110010010001111110000,
32'b 00000011110110111010011000010000,
32'b 00011111011110111010101001100000,
32'b 00000011000111101111001110000000,
32'b 00011111000111000110001011110000,
32'b 00000000000000000000000000000000,
32'b 00000000000000011000000000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000111111111100000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000000111100000000000000,
32'b 00000000000011111110001111000000,
32'b 00000000000011111110111101000000,
32'b 00000000000111111111111011100000,
32'b 00000000000111111111110111110000,
32'b 00000000001111111111110011100000,
32'b 00000000001111111111010001000000,
32'b 00000000000111111111010000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000001111110000000000000,
32'b 00000000000001111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000001111111111100000000000,


32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00011111001110010010001111110000,
32'b 00000011110110111010011000010000,
32'b 00011111011110111010101001100000,
32'b 00000011000111101111001110000000,
32'b 00011111000111000110001011110000,
32'b 00000000000000000000000000000000,
32'b 00000000000000011000000000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000111111111100000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000000111100000000000000,
32'b 00000000000011111110001111000000,
32'b 00000000000011111110111101000000,
32'b 00000000000111111111111011100000,
32'b 00000000000111111111110111110000,
32'b 00000000001111111111110011100000,
32'b 00000000001111111111010001000000,
32'b 00000000000111111111010000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000001111110000000000000,
32'b 00000000000001111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000001111111111100000000000,
		
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00011111001110010010001111110000,
32'b 00000011110110111010011000010000,
32'b 00011111011110111010101001100000,
32'b 00000011000111101111001110000000,
32'b 00011111000111000110001011110000,
32'b 00000000000000000000000000000000,
32'b 00000000000000011000000000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000111111111100000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000000111100000000000000,
32'b 00000000000011111110001111000000,
32'b 00000000000011111110111101000000,
32'b 00000000000111111111111011100000,
32'b 00000000000111111111110111110000,
32'b 00000000001111111111110011100000,
32'b 00000000001111111111010001000000,
32'b 00000000000111111111010000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000001111110000000000000,
32'b 00000000000001111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000001111111111100000000000,
		
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00000000000000000000000000000000,
32'b 00011111001110010010001111110000,
32'b 00000011110110111010011000010000,
32'b 00011111011110111010101001100000,
32'b 00000011000111101111001110000000,
32'b 00011111000111000110001011110000,
32'b 00000000000000000000000000000000,
32'b 00000000000000011000000000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000111111111100000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000000111100000000000000,
32'b 00000000000011111110001111000000,
32'b 00000000000011111110111101000000,
32'b 00000000000111111111111011100000,
32'b 00000000000111111111110111110000,
32'b 00000000001111111111110011100000,
32'b 00000000001111111111010001000000,
32'b 00000000000111111111010000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000011111111000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000000001111110000000000000,
32'b 00000000000001111110000000000000,
32'b 00000000000011111110000000000000,
32'b 00000000001111111111100000000000
		


	};

	assign data = ROM[addr];

endmodule
